** Profile: "SCHEMATIC1-pwmSmoothingTest"  [ D:\DROPBOX\CLASSES\ME 344\Maglev lab - Group Files\pwmToAnalogConverter-PSpiceFiles\SCHEMATIC1\pwmSmoothingTest.sim ] 

** Creating circuit file "pwmSmoothingTest.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\Justin\AppData\Roaming\SPB_16.6\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 0.1s 0 500ns 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
